module main

struct Data_control {
	state i8
	mod_by string
	created_by string
}
